`include "types.sv"

